magic
tech sky130A
magscale 1 2
timestamp 1695510773
<< viali >>
rect 2237 7905 2271 7939
rect 2789 7837 2823 7871
rect 6193 7837 6227 7871
rect 6653 7837 6687 7871
rect 6469 7769 6503 7803
rect 4248 6953 4282 6987
rect 5733 6817 5767 6851
rect 2881 6749 2915 6783
rect 3341 6749 3375 6783
rect 3985 6749 4019 6783
rect 2614 6681 2648 6715
rect 1501 6613 1535 6647
rect 3249 6613 3283 6647
rect 4077 6409 4111 6443
rect 5733 6409 5767 6443
rect 5365 6341 5399 6375
rect 2789 6273 2823 6307
rect 5089 6273 5123 6307
rect 5825 6273 5859 6307
rect 4905 6205 4939 6239
rect 4997 6205 5031 6239
rect 5181 6205 5215 6239
rect 3525 5865 3559 5899
rect 3893 5797 3927 5831
rect 2053 5729 2087 5763
rect 1777 5661 1811 5695
rect 4077 5661 4111 5695
rect 4077 5321 4111 5355
rect 2513 5185 2547 5219
rect 2789 5185 2823 5219
rect 2421 4981 2455 5015
rect 5549 4777 5583 4811
rect 4905 4641 4939 4675
rect 4077 4573 4111 4607
rect 4261 4573 4295 4607
rect 4353 4573 4387 4607
rect 4629 4573 4663 4607
rect 4721 4573 4755 4607
rect 5457 4573 5491 4607
rect 5641 4573 5675 4607
rect 5917 4573 5951 4607
rect 6101 4573 6135 4607
rect 2605 4437 2639 4471
rect 3893 4437 3927 4471
rect 4905 4437 4939 4471
rect 6009 4437 6043 4471
rect 3801 4233 3835 4267
rect 1501 4097 1535 4131
rect 3893 4097 3927 4131
rect 4629 4097 4663 4131
rect 5181 4097 5215 4131
rect 5641 4097 5675 4131
rect 5825 4097 5859 4131
rect 1777 4029 1811 4063
rect 3709 4029 3743 4063
rect 4813 4029 4847 4063
rect 4905 4029 4939 4063
rect 5457 4029 5491 4063
rect 5917 4029 5951 4063
rect 4261 3961 4295 3995
rect 4721 3961 4755 3995
rect 3249 3893 3283 3927
rect 4997 3893 5031 3927
rect 3525 3689 3559 3723
rect 4997 3689 5031 3723
rect 3433 3621 3467 3655
rect 3065 3553 3099 3587
rect 5641 3553 5675 3587
rect 3985 3485 4019 3519
rect 5457 3417 5491 3451
rect 4077 3349 4111 3383
rect 5365 3349 5399 3383
rect 1777 3145 1811 3179
rect 4537 3145 4571 3179
rect 3249 3077 3283 3111
rect 3801 3077 3835 3111
rect 3985 3009 4019 3043
rect 4077 3009 4111 3043
rect 4445 3009 4479 3043
rect 4629 3009 4663 3043
rect 3801 2873 3835 2907
rect 5825 2465 5859 2499
rect 6101 2397 6135 2431
rect 6653 2261 6687 2295
<< metal1 >>
rect 1104 8186 7176 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 7176 8186
rect 1104 8112 7176 8134
rect 2774 8072 2780 8084
rect 2746 8032 2780 8072
rect 2832 8032 2838 8084
rect 2225 7939 2283 7945
rect 2225 7905 2237 7939
rect 2271 7936 2283 7939
rect 2746 7936 2774 8032
rect 2271 7908 2774 7936
rect 2271 7905 2283 7908
rect 2225 7899 2283 7905
rect 2774 7828 2780 7880
rect 2832 7828 2838 7880
rect 6181 7871 6239 7877
rect 6181 7837 6193 7871
rect 6227 7868 6239 7871
rect 6641 7871 6699 7877
rect 6641 7868 6653 7871
rect 6227 7840 6653 7868
rect 6227 7837 6239 7840
rect 6181 7831 6239 7837
rect 6641 7837 6653 7840
rect 6687 7868 6699 7871
rect 7742 7868 7748 7880
rect 6687 7840 7748 7868
rect 6687 7837 6699 7840
rect 6641 7831 6699 7837
rect 7742 7828 7748 7840
rect 7800 7828 7806 7880
rect 6454 7760 6460 7812
rect 6512 7760 6518 7812
rect 1104 7642 7176 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 7176 7642
rect 1104 7568 7176 7590
rect 1104 7098 7176 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 7176 7098
rect 1104 7024 7176 7046
rect 4236 6987 4294 6993
rect 4236 6953 4248 6987
rect 4282 6984 4294 6987
rect 4706 6984 4712 6996
rect 4282 6956 4712 6984
rect 4282 6953 4294 6956
rect 4236 6947 4294 6953
rect 4706 6944 4712 6956
rect 4764 6944 4770 6996
rect 4798 6808 4804 6860
rect 4856 6848 4862 6860
rect 5721 6851 5779 6857
rect 5721 6848 5733 6851
rect 4856 6820 5733 6848
rect 4856 6808 4862 6820
rect 5721 6817 5733 6820
rect 5767 6817 5779 6851
rect 5721 6811 5779 6817
rect 2869 6783 2927 6789
rect 2869 6749 2881 6783
rect 2915 6749 2927 6783
rect 2869 6743 2927 6749
rect 3329 6783 3387 6789
rect 3329 6749 3341 6783
rect 3375 6780 3387 6783
rect 3878 6780 3884 6792
rect 3375 6752 3884 6780
rect 3375 6749 3387 6752
rect 3329 6743 3387 6749
rect 2590 6672 2596 6724
rect 2648 6721 2654 6724
rect 2648 6675 2660 6721
rect 2884 6712 2912 6743
rect 3878 6740 3884 6752
rect 3936 6740 3942 6792
rect 3973 6783 4031 6789
rect 3973 6749 3985 6783
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 3988 6712 4016 6743
rect 5534 6712 5540 6724
rect 2884 6684 4108 6712
rect 5474 6684 5540 6712
rect 2648 6672 2654 6675
rect 4080 6656 4108 6684
rect 5534 6672 5540 6684
rect 5592 6672 5598 6724
rect 1489 6647 1547 6653
rect 1489 6613 1501 6647
rect 1535 6644 1547 6647
rect 2774 6644 2780 6656
rect 1535 6616 2780 6644
rect 1535 6613 1547 6616
rect 1489 6607 1547 6613
rect 2774 6604 2780 6616
rect 2832 6604 2838 6656
rect 3142 6604 3148 6656
rect 3200 6644 3206 6656
rect 3237 6647 3295 6653
rect 3237 6644 3249 6647
rect 3200 6616 3249 6644
rect 3200 6604 3206 6616
rect 3237 6613 3249 6616
rect 3283 6613 3295 6647
rect 3237 6607 3295 6613
rect 4062 6604 4068 6656
rect 4120 6604 4126 6656
rect 1104 6554 7176 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 7176 6554
rect 1104 6480 7176 6502
rect 2590 6400 2596 6452
rect 2648 6400 2654 6452
rect 4062 6400 4068 6452
rect 4120 6400 4126 6452
rect 5534 6400 5540 6452
rect 5592 6440 5598 6452
rect 5721 6443 5779 6449
rect 5721 6440 5733 6443
rect 5592 6412 5733 6440
rect 5592 6400 5598 6412
rect 5721 6409 5733 6412
rect 5767 6409 5779 6443
rect 5721 6403 5779 6409
rect 6454 6400 6460 6452
rect 6512 6400 6518 6452
rect 2608 6372 2636 6400
rect 5353 6375 5411 6381
rect 5353 6372 5365 6375
rect 2608 6344 5365 6372
rect 5353 6341 5365 6344
rect 5399 6341 5411 6375
rect 5353 6335 5411 6341
rect 2774 6264 2780 6316
rect 2832 6264 2838 6316
rect 3878 6264 3884 6316
rect 3936 6304 3942 6316
rect 5077 6307 5135 6313
rect 5077 6304 5089 6307
rect 3936 6276 5089 6304
rect 3936 6264 3942 6276
rect 5077 6273 5089 6276
rect 5123 6304 5135 6307
rect 5813 6307 5871 6313
rect 5813 6304 5825 6307
rect 5123 6276 5825 6304
rect 5123 6273 5135 6276
rect 5077 6267 5135 6273
rect 5813 6273 5825 6276
rect 5859 6304 5871 6307
rect 6472 6304 6500 6400
rect 5859 6276 6500 6304
rect 5859 6273 5871 6276
rect 5813 6267 5871 6273
rect 4798 6196 4804 6248
rect 4856 6236 4862 6248
rect 4893 6239 4951 6245
rect 4893 6236 4905 6239
rect 4856 6208 4905 6236
rect 4856 6196 4862 6208
rect 4893 6205 4905 6208
rect 4939 6205 4951 6239
rect 4893 6199 4951 6205
rect 4985 6239 5043 6245
rect 4985 6205 4997 6239
rect 5031 6205 5043 6239
rect 4985 6199 5043 6205
rect 5169 6239 5227 6245
rect 5169 6205 5181 6239
rect 5215 6236 5227 6239
rect 5534 6236 5540 6248
rect 5215 6208 5540 6236
rect 5215 6205 5227 6208
rect 5169 6199 5227 6205
rect 3510 6128 3516 6180
rect 3568 6168 3574 6180
rect 5000 6168 5028 6199
rect 5534 6196 5540 6208
rect 5592 6196 5598 6248
rect 3568 6140 5028 6168
rect 3568 6128 3574 6140
rect 1104 6010 7176 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 7176 6010
rect 1104 5936 7176 5958
rect 3510 5856 3516 5908
rect 3568 5856 3574 5908
rect 3881 5831 3939 5837
rect 3881 5797 3893 5831
rect 3927 5797 3939 5831
rect 3881 5791 3939 5797
rect 2041 5763 2099 5769
rect 2041 5729 2053 5763
rect 2087 5760 2099 5763
rect 3896 5760 3924 5791
rect 2087 5732 3924 5760
rect 2087 5729 2099 5732
rect 2041 5723 2099 5729
rect 1486 5652 1492 5704
rect 1544 5692 1550 5704
rect 1765 5695 1823 5701
rect 1765 5692 1777 5695
rect 1544 5664 1777 5692
rect 1544 5652 1550 5664
rect 1765 5661 1777 5664
rect 1811 5661 1823 5695
rect 1765 5655 1823 5661
rect 3142 5652 3148 5704
rect 3200 5652 3206 5704
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5692 4123 5695
rect 4614 5692 4620 5704
rect 4111 5664 4620 5692
rect 4111 5661 4123 5664
rect 4065 5655 4123 5661
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 1104 5466 7176 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 7176 5466
rect 1104 5392 7176 5414
rect 2774 5312 2780 5364
rect 2832 5352 2838 5364
rect 3234 5352 3240 5364
rect 2832 5324 3240 5352
rect 2832 5312 2838 5324
rect 3234 5312 3240 5324
rect 3292 5352 3298 5364
rect 4065 5355 4123 5361
rect 4065 5352 4077 5355
rect 3292 5324 4077 5352
rect 3292 5312 3298 5324
rect 4065 5321 4077 5324
rect 4111 5321 4123 5355
rect 4065 5315 4123 5321
rect 3878 5284 3884 5296
rect 2516 5256 3884 5284
rect 2516 5225 2544 5256
rect 3878 5244 3884 5256
rect 3936 5244 3942 5296
rect 2501 5219 2559 5225
rect 2501 5185 2513 5219
rect 2547 5185 2559 5219
rect 2777 5219 2835 5225
rect 2777 5216 2789 5219
rect 2501 5179 2559 5185
rect 2608 5188 2789 5216
rect 2608 5024 2636 5188
rect 2777 5185 2789 5188
rect 2823 5185 2835 5219
rect 2777 5179 2835 5185
rect 2406 4972 2412 5024
rect 2464 4972 2470 5024
rect 2590 4972 2596 5024
rect 2648 4972 2654 5024
rect 1104 4922 7176 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 7176 4922
rect 1104 4848 7176 4870
rect 5258 4768 5264 4820
rect 5316 4808 5322 4820
rect 5316 4780 5488 4808
rect 5316 4768 5322 4780
rect 5350 4740 5356 4752
rect 4816 4712 5356 4740
rect 4816 4684 4844 4712
rect 5350 4700 5356 4712
rect 5408 4700 5414 4752
rect 5460 4740 5488 4780
rect 5534 4768 5540 4820
rect 5592 4768 5598 4820
rect 5460 4712 5948 4740
rect 4798 4672 4804 4684
rect 4632 4644 4804 4672
rect 4065 4607 4123 4613
rect 4065 4573 4077 4607
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 4080 4536 4108 4567
rect 4246 4564 4252 4616
rect 4304 4564 4310 4616
rect 4338 4564 4344 4616
rect 4396 4564 4402 4616
rect 4632 4613 4660 4644
rect 4798 4632 4804 4644
rect 4856 4632 4862 4684
rect 4893 4675 4951 4681
rect 4893 4641 4905 4675
rect 4939 4672 4951 4675
rect 5166 4672 5172 4684
rect 4939 4644 5172 4672
rect 4939 4641 4951 4644
rect 4893 4635 4951 4641
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 4617 4607 4675 4613
rect 4617 4573 4629 4607
rect 4663 4573 4675 4607
rect 4617 4567 4675 4573
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4604 4767 4607
rect 5258 4604 5264 4616
rect 4755 4576 5264 4604
rect 4755 4573 4767 4576
rect 4709 4567 4767 4573
rect 5258 4564 5264 4576
rect 5316 4604 5322 4616
rect 5920 4613 5948 4712
rect 5445 4607 5503 4613
rect 5445 4604 5457 4607
rect 5316 4576 5457 4604
rect 5316 4564 5322 4576
rect 5445 4573 5457 4576
rect 5491 4573 5503 4607
rect 5445 4567 5503 4573
rect 5629 4607 5687 4613
rect 5629 4573 5641 4607
rect 5675 4604 5687 4607
rect 5905 4607 5963 4613
rect 5675 4576 5764 4604
rect 5675 4573 5687 4576
rect 5629 4567 5687 4573
rect 4798 4536 4804 4548
rect 4080 4508 4804 4536
rect 4798 4496 4804 4508
rect 4856 4496 4862 4548
rect 5736 4536 5764 4576
rect 5905 4573 5917 4607
rect 5951 4573 5963 4607
rect 5905 4567 5963 4573
rect 6089 4607 6147 4613
rect 6089 4573 6101 4607
rect 6135 4573 6147 4607
rect 6089 4567 6147 4573
rect 6104 4536 6132 4567
rect 5736 4508 6132 4536
rect 5736 4480 5764 4508
rect 14 4428 20 4480
rect 72 4468 78 4480
rect 2590 4468 2596 4480
rect 72 4440 2596 4468
rect 72 4428 78 4440
rect 2590 4428 2596 4440
rect 2648 4428 2654 4480
rect 3326 4428 3332 4480
rect 3384 4468 3390 4480
rect 3881 4471 3939 4477
rect 3881 4468 3893 4471
rect 3384 4440 3893 4468
rect 3384 4428 3390 4440
rect 3881 4437 3893 4440
rect 3927 4437 3939 4471
rect 3881 4431 3939 4437
rect 4154 4428 4160 4480
rect 4212 4468 4218 4480
rect 4893 4471 4951 4477
rect 4893 4468 4905 4471
rect 4212 4440 4905 4468
rect 4212 4428 4218 4440
rect 4893 4437 4905 4440
rect 4939 4437 4951 4471
rect 4893 4431 4951 4437
rect 5166 4428 5172 4480
rect 5224 4468 5230 4480
rect 5718 4468 5724 4480
rect 5224 4440 5724 4468
rect 5224 4428 5230 4440
rect 5718 4428 5724 4440
rect 5776 4428 5782 4480
rect 5994 4428 6000 4480
rect 6052 4428 6058 4480
rect 1104 4378 7176 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 7176 4378
rect 1104 4304 7176 4326
rect 3786 4224 3792 4276
rect 3844 4264 3850 4276
rect 4246 4264 4252 4276
rect 3844 4236 4252 4264
rect 3844 4224 3850 4236
rect 4246 4224 4252 4236
rect 4304 4224 4310 4276
rect 2406 4156 2412 4208
rect 2464 4156 2470 4208
rect 5184 4168 5764 4196
rect 1486 4088 1492 4140
rect 1544 4088 1550 4140
rect 3510 4088 3516 4140
rect 3568 4128 3574 4140
rect 3568 4100 3832 4128
rect 3568 4088 3574 4100
rect 1765 4063 1823 4069
rect 1765 4029 1777 4063
rect 1811 4060 1823 4063
rect 3326 4060 3332 4072
rect 1811 4032 3332 4060
rect 1811 4029 1823 4032
rect 1765 4023 1823 4029
rect 3326 4020 3332 4032
rect 3384 4020 3390 4072
rect 3697 4063 3755 4069
rect 3697 4029 3709 4063
rect 3743 4029 3755 4063
rect 3804 4060 3832 4100
rect 3878 4088 3884 4140
rect 3936 4088 3942 4140
rect 5184 4137 5212 4168
rect 5736 4140 5764 4168
rect 4617 4131 4675 4137
rect 4080 4100 4292 4128
rect 4080 4060 4108 4100
rect 3804 4032 4108 4060
rect 3697 4023 3755 4029
rect 3712 3992 3740 4023
rect 4154 4020 4160 4072
rect 4212 4020 4218 4072
rect 4264 4060 4292 4100
rect 4617 4097 4629 4131
rect 4663 4128 4675 4131
rect 5169 4131 5227 4137
rect 4663 4100 5028 4128
rect 4663 4097 4675 4100
rect 4617 4091 4675 4097
rect 4801 4063 4859 4069
rect 4801 4060 4813 4063
rect 4264 4032 4813 4060
rect 4801 4029 4813 4032
rect 4847 4029 4859 4063
rect 4801 4023 4859 4029
rect 4893 4063 4951 4069
rect 4893 4029 4905 4063
rect 4939 4029 4951 4063
rect 5000 4060 5028 4100
rect 5169 4097 5181 4131
rect 5215 4097 5227 4131
rect 5169 4091 5227 4097
rect 5534 4088 5540 4140
rect 5592 4128 5598 4140
rect 5629 4131 5687 4137
rect 5629 4128 5641 4131
rect 5592 4100 5641 4128
rect 5592 4088 5598 4100
rect 5629 4097 5641 4100
rect 5675 4097 5687 4131
rect 5629 4091 5687 4097
rect 5718 4088 5724 4140
rect 5776 4088 5782 4140
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 5994 4128 6000 4140
rect 5859 4100 6000 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 5994 4088 6000 4100
rect 6052 4088 6058 4140
rect 5445 4063 5503 4069
rect 5445 4060 5457 4063
rect 5000 4032 5457 4060
rect 4893 4023 4951 4029
rect 5445 4029 5457 4032
rect 5491 4029 5503 4063
rect 5445 4023 5503 4029
rect 5905 4063 5963 4069
rect 5905 4029 5917 4063
rect 5951 4029 5963 4063
rect 5905 4023 5963 4029
rect 4172 3992 4200 4020
rect 3712 3964 4200 3992
rect 4249 3995 4307 4001
rect 4249 3961 4261 3995
rect 4295 3992 4307 3995
rect 4614 3992 4620 4004
rect 4295 3964 4620 3992
rect 4295 3961 4307 3964
rect 4249 3955 4307 3961
rect 4614 3952 4620 3964
rect 4672 3952 4678 4004
rect 4706 3952 4712 4004
rect 4764 3952 4770 4004
rect 3050 3884 3056 3936
rect 3108 3924 3114 3936
rect 3237 3927 3295 3933
rect 3237 3924 3249 3927
rect 3108 3896 3249 3924
rect 3108 3884 3114 3896
rect 3237 3893 3249 3896
rect 3283 3893 3295 3927
rect 3237 3887 3295 3893
rect 4338 3884 4344 3936
rect 4396 3924 4402 3936
rect 4798 3924 4804 3936
rect 4396 3896 4804 3924
rect 4396 3884 4402 3896
rect 4798 3884 4804 3896
rect 4856 3924 4862 3936
rect 4908 3924 4936 4023
rect 5350 3952 5356 4004
rect 5408 3992 5414 4004
rect 5920 3992 5948 4023
rect 5408 3964 5948 3992
rect 5408 3952 5414 3964
rect 4856 3896 4936 3924
rect 4856 3884 4862 3896
rect 4982 3884 4988 3936
rect 5040 3924 5046 3936
rect 5258 3924 5264 3936
rect 5040 3896 5264 3924
rect 5040 3884 5046 3896
rect 5258 3884 5264 3896
rect 5316 3884 5322 3936
rect 1104 3834 7176 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 7176 3834
rect 1104 3760 7176 3782
rect 3050 3680 3056 3732
rect 3108 3680 3114 3732
rect 3513 3723 3571 3729
rect 3513 3689 3525 3723
rect 3559 3720 3571 3723
rect 3786 3720 3792 3732
rect 3559 3692 3792 3720
rect 3559 3689 3571 3692
rect 3513 3683 3571 3689
rect 3786 3680 3792 3692
rect 3844 3680 3850 3732
rect 4890 3680 4896 3732
rect 4948 3720 4954 3732
rect 4985 3723 5043 3729
rect 4985 3720 4997 3723
rect 4948 3692 4997 3720
rect 4948 3680 4954 3692
rect 4985 3689 4997 3692
rect 5031 3689 5043 3723
rect 4985 3683 5043 3689
rect 3068 3593 3096 3680
rect 3418 3612 3424 3664
rect 3476 3612 3482 3664
rect 3053 3587 3111 3593
rect 3053 3553 3065 3587
rect 3099 3584 3111 3587
rect 3099 3556 4016 3584
rect 3099 3553 3111 3556
rect 3053 3547 3111 3553
rect 3988 3525 4016 3556
rect 5350 3544 5356 3596
rect 5408 3544 5414 3596
rect 5629 3587 5687 3593
rect 5629 3553 5641 3587
rect 5675 3584 5687 3587
rect 5810 3584 5816 3596
rect 5675 3556 5816 3584
rect 5675 3553 5687 3556
rect 5629 3547 5687 3553
rect 5810 3544 5816 3556
rect 5868 3544 5874 3596
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 5368 3448 5396 3544
rect 5445 3451 5503 3457
rect 5445 3448 5457 3451
rect 5368 3420 5457 3448
rect 5445 3417 5457 3420
rect 5491 3417 5503 3451
rect 5445 3411 5503 3417
rect 4062 3340 4068 3392
rect 4120 3380 4126 3392
rect 4982 3380 4988 3392
rect 4120 3352 4988 3380
rect 4120 3340 4126 3352
rect 4982 3340 4988 3352
rect 5040 3380 5046 3392
rect 5353 3383 5411 3389
rect 5353 3380 5365 3383
rect 5040 3352 5365 3380
rect 5040 3340 5046 3352
rect 5353 3349 5365 3352
rect 5399 3349 5411 3383
rect 5353 3343 5411 3349
rect 1104 3290 7176 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 7176 3290
rect 1104 3216 7176 3238
rect 1486 3136 1492 3188
rect 1544 3176 1550 3188
rect 1765 3179 1823 3185
rect 1765 3176 1777 3179
rect 1544 3148 1777 3176
rect 1544 3136 1550 3148
rect 1765 3145 1777 3148
rect 1811 3145 1823 3179
rect 1765 3139 1823 3145
rect 4525 3179 4583 3185
rect 4525 3145 4537 3179
rect 4571 3176 4583 3179
rect 4798 3176 4804 3188
rect 4571 3148 4804 3176
rect 4571 3145 4583 3148
rect 4525 3139 4583 3145
rect 4798 3136 4804 3148
rect 4856 3136 4862 3188
rect 3234 3068 3240 3120
rect 3292 3068 3298 3120
rect 3418 3068 3424 3120
rect 3476 3108 3482 3120
rect 3789 3111 3847 3117
rect 3789 3108 3801 3111
rect 3476 3080 3801 3108
rect 3476 3068 3482 3080
rect 3789 3077 3801 3080
rect 3835 3108 3847 3111
rect 3835 3080 4476 3108
rect 3835 3077 3847 3080
rect 3789 3071 3847 3077
rect 3973 3043 4031 3049
rect 3973 3009 3985 3043
rect 4019 3009 4031 3043
rect 3973 3003 4031 3009
rect 3878 2932 3884 2984
rect 3936 2932 3942 2984
rect 3988 2972 4016 3003
rect 4062 3000 4068 3052
rect 4120 3000 4126 3052
rect 4448 3049 4476 3080
rect 4433 3043 4491 3049
rect 4433 3009 4445 3043
rect 4479 3009 4491 3043
rect 4433 3003 4491 3009
rect 4617 3043 4675 3049
rect 4617 3009 4629 3043
rect 4663 3040 4675 3043
rect 5350 3040 5356 3052
rect 4663 3012 5356 3040
rect 4663 3009 4675 3012
rect 4617 3003 4675 3009
rect 4632 2972 4660 3003
rect 5350 3000 5356 3012
rect 5408 3000 5414 3052
rect 3988 2944 4660 2972
rect 3789 2907 3847 2913
rect 3789 2873 3801 2907
rect 3835 2904 3847 2907
rect 3896 2904 3924 2932
rect 3835 2876 3924 2904
rect 3835 2873 3847 2876
rect 3789 2867 3847 2873
rect 1104 2746 7176 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 7176 2746
rect 1104 2672 7176 2694
rect 5810 2456 5816 2508
rect 5868 2456 5874 2508
rect 6089 2431 6147 2437
rect 6089 2397 6101 2431
rect 6135 2428 6147 2431
rect 6135 2400 6684 2428
rect 6135 2397 6147 2400
rect 6089 2391 6147 2397
rect 6656 2304 6684 2400
rect 6638 2252 6644 2304
rect 6696 2252 6702 2304
rect 1104 2202 7176 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 7176 2202
rect 1104 2128 7176 2150
<< via1 >>
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 2780 8032 2832 8084
rect 2780 7871 2832 7880
rect 2780 7837 2789 7871
rect 2789 7837 2823 7871
rect 2823 7837 2832 7871
rect 2780 7828 2832 7837
rect 7748 7828 7800 7880
rect 6460 7803 6512 7812
rect 6460 7769 6469 7803
rect 6469 7769 6503 7803
rect 6503 7769 6512 7803
rect 6460 7760 6512 7769
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 4712 6944 4764 6996
rect 4804 6808 4856 6860
rect 2596 6715 2648 6724
rect 2596 6681 2614 6715
rect 2614 6681 2648 6715
rect 2596 6672 2648 6681
rect 3884 6740 3936 6792
rect 5540 6672 5592 6724
rect 2780 6604 2832 6656
rect 3148 6604 3200 6656
rect 4068 6604 4120 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 2596 6400 2648 6452
rect 4068 6443 4120 6452
rect 4068 6409 4077 6443
rect 4077 6409 4111 6443
rect 4111 6409 4120 6443
rect 4068 6400 4120 6409
rect 5540 6400 5592 6452
rect 6460 6400 6512 6452
rect 2780 6307 2832 6316
rect 2780 6273 2789 6307
rect 2789 6273 2823 6307
rect 2823 6273 2832 6307
rect 2780 6264 2832 6273
rect 3884 6264 3936 6316
rect 4804 6196 4856 6248
rect 3516 6128 3568 6180
rect 5540 6196 5592 6248
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 3516 5899 3568 5908
rect 3516 5865 3525 5899
rect 3525 5865 3559 5899
rect 3559 5865 3568 5899
rect 3516 5856 3568 5865
rect 1492 5652 1544 5704
rect 3148 5652 3200 5704
rect 4620 5652 4672 5704
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 2780 5312 2832 5364
rect 3240 5312 3292 5364
rect 3884 5244 3936 5296
rect 2412 5015 2464 5024
rect 2412 4981 2421 5015
rect 2421 4981 2455 5015
rect 2455 4981 2464 5015
rect 2412 4972 2464 4981
rect 2596 4972 2648 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 5264 4768 5316 4820
rect 5356 4700 5408 4752
rect 5540 4811 5592 4820
rect 5540 4777 5549 4811
rect 5549 4777 5583 4811
rect 5583 4777 5592 4811
rect 5540 4768 5592 4777
rect 4252 4607 4304 4616
rect 4252 4573 4261 4607
rect 4261 4573 4295 4607
rect 4295 4573 4304 4607
rect 4252 4564 4304 4573
rect 4344 4607 4396 4616
rect 4344 4573 4353 4607
rect 4353 4573 4387 4607
rect 4387 4573 4396 4607
rect 4344 4564 4396 4573
rect 4804 4632 4856 4684
rect 5172 4632 5224 4684
rect 5264 4564 5316 4616
rect 4804 4496 4856 4548
rect 20 4428 72 4480
rect 2596 4471 2648 4480
rect 2596 4437 2605 4471
rect 2605 4437 2639 4471
rect 2639 4437 2648 4471
rect 2596 4428 2648 4437
rect 3332 4428 3384 4480
rect 4160 4428 4212 4480
rect 5172 4428 5224 4480
rect 5724 4428 5776 4480
rect 6000 4471 6052 4480
rect 6000 4437 6009 4471
rect 6009 4437 6043 4471
rect 6043 4437 6052 4471
rect 6000 4428 6052 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 3792 4267 3844 4276
rect 3792 4233 3801 4267
rect 3801 4233 3835 4267
rect 3835 4233 3844 4267
rect 3792 4224 3844 4233
rect 4252 4224 4304 4276
rect 2412 4156 2464 4208
rect 1492 4131 1544 4140
rect 1492 4097 1501 4131
rect 1501 4097 1535 4131
rect 1535 4097 1544 4131
rect 1492 4088 1544 4097
rect 3516 4088 3568 4140
rect 3332 4020 3384 4072
rect 3884 4131 3936 4140
rect 3884 4097 3893 4131
rect 3893 4097 3927 4131
rect 3927 4097 3936 4131
rect 3884 4088 3936 4097
rect 4160 4020 4212 4072
rect 5540 4088 5592 4140
rect 5724 4088 5776 4140
rect 6000 4088 6052 4140
rect 4620 3952 4672 4004
rect 4712 3995 4764 4004
rect 4712 3961 4721 3995
rect 4721 3961 4755 3995
rect 4755 3961 4764 3995
rect 4712 3952 4764 3961
rect 3056 3884 3108 3936
rect 4344 3884 4396 3936
rect 4804 3884 4856 3936
rect 5356 3952 5408 4004
rect 4988 3927 5040 3936
rect 4988 3893 4997 3927
rect 4997 3893 5031 3927
rect 5031 3893 5040 3927
rect 4988 3884 5040 3893
rect 5264 3884 5316 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 3056 3680 3108 3732
rect 3792 3680 3844 3732
rect 4896 3680 4948 3732
rect 3424 3655 3476 3664
rect 3424 3621 3433 3655
rect 3433 3621 3467 3655
rect 3467 3621 3476 3655
rect 3424 3612 3476 3621
rect 5356 3544 5408 3596
rect 5816 3544 5868 3596
rect 4068 3383 4120 3392
rect 4068 3349 4077 3383
rect 4077 3349 4111 3383
rect 4111 3349 4120 3383
rect 4068 3340 4120 3349
rect 4988 3340 5040 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 1492 3136 1544 3188
rect 4804 3136 4856 3188
rect 3240 3111 3292 3120
rect 3240 3077 3249 3111
rect 3249 3077 3283 3111
rect 3283 3077 3292 3111
rect 3240 3068 3292 3077
rect 3424 3068 3476 3120
rect 3884 2932 3936 2984
rect 4068 3043 4120 3052
rect 4068 3009 4077 3043
rect 4077 3009 4111 3043
rect 4111 3009 4120 3043
rect 4068 3000 4120 3009
rect 5356 3000 5408 3052
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 5816 2499 5868 2508
rect 5816 2465 5825 2499
rect 5825 2465 5859 2499
rect 5859 2465 5868 2499
rect 5816 2456 5868 2465
rect 6644 2295 6696 2304
rect 6644 2261 6653 2295
rect 6653 2261 6687 2295
rect 6687 2261 6696 2295
rect 6644 2252 6696 2261
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 7746 9687 7802 10487
rect 2778 9616 2834 9625
rect 2778 9551 2834 9560
rect 2792 8090 2820 9551
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 7760 7886 7788 9687
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 2596 6724 2648 6730
rect 2596 6666 2648 6672
rect 2608 6458 2636 6666
rect 2792 6662 2820 7822
rect 6460 7812 6512 7818
rect 6460 7754 6512 7760
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4712 6996 4764 7002
rect 4712 6938 4764 6944
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 1492 5704 1544 5710
rect 1492 5646 1544 5652
rect 20 4480 72 4486
rect 20 4422 72 4428
rect 32 800 60 4422
rect 1504 4146 1532 5646
rect 2792 5370 2820 6258
rect 3160 5710 3188 6598
rect 3896 6322 3924 6734
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 4080 6458 4108 6598
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 3516 6180 3568 6186
rect 3516 6122 3568 6128
rect 3528 5914 3556 6122
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 2412 5024 2464 5030
rect 2412 4966 2464 4972
rect 2596 5024 2648 5030
rect 2596 4966 2648 4972
rect 2424 4214 2452 4966
rect 2608 4486 2636 4966
rect 2596 4480 2648 4486
rect 2596 4422 2648 4428
rect 2412 4208 2464 4214
rect 2412 4150 2464 4156
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1504 3194 1532 4082
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 3068 3738 3096 3878
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 1492 3188 1544 3194
rect 1492 3130 1544 3136
rect 3252 3126 3280 5306
rect 3332 4480 3384 4486
rect 3332 4422 3384 4428
rect 3344 4078 3372 4422
rect 3528 4146 3556 5850
rect 3896 5302 3924 6258
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 3792 4276 3844 4282
rect 3792 4218 3844 4224
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 3332 4072 3384 4078
rect 3528 4026 3556 4082
rect 3332 4014 3384 4020
rect 3436 3998 3556 4026
rect 3436 3670 3464 3998
rect 3804 3738 3832 4218
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3424 3664 3476 3670
rect 3424 3606 3476 3612
rect 3436 3126 3464 3606
rect 3240 3120 3292 3126
rect 3240 3062 3292 3068
rect 3424 3120 3476 3126
rect 3424 3062 3476 3068
rect 3896 2990 3924 4082
rect 4172 4078 4200 4422
rect 4264 4282 4292 4558
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 4356 3942 4384 4558
rect 4632 4010 4660 5646
rect 4724 4010 4752 6938
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4816 6254 4844 6802
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 5552 6458 5580 6666
rect 6472 6458 6500 7754
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 4816 4690 4844 6190
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 5552 4826 5580 6190
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 4804 4548 4856 4554
rect 4804 4490 4856 4496
rect 4816 4026 4844 4490
rect 5184 4486 5212 4626
rect 5276 4622 5304 4762
rect 5356 4752 5408 4758
rect 5356 4694 5408 4700
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4712 4004 4764 4010
rect 4816 3998 4936 4026
rect 4712 3946 4764 3952
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 4080 3058 4108 3334
rect 4816 3194 4844 3878
rect 4908 3738 4936 3998
rect 5276 3942 5304 4558
rect 5368 4010 5396 4694
rect 5552 4146 5580 4762
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 5736 4146 5764 4422
rect 6012 4146 6040 4422
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5724 4140 5776 4146
rect 6000 4140 6052 4146
rect 5776 4100 5856 4128
rect 5724 4082 5776 4088
rect 5356 4004 5408 4010
rect 5356 3946 5408 3952
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 5000 3398 5028 3878
rect 5368 3602 5396 3946
rect 5828 3602 5856 4100
rect 6000 4082 6052 4088
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 5816 3596 5868 3602
rect 5816 3538 5868 3544
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 5368 3058 5396 3538
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 3884 2984 3936 2990
rect 3884 2926 3936 2932
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 5828 2514 5856 3538
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 6644 2304 6696 2310
rect 6644 2246 6696 2252
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 18 0 74 800
rect 6656 785 6684 2246
rect 6642 776 6698 785
rect 6642 711 6698 720
<< via2 >>
rect 2778 9560 2834 9616
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 6642 720 6698 776
<< metal3 >>
rect 0 9618 800 9648
rect 2773 9618 2839 9621
rect 0 9616 2839 9618
rect 0 9560 2778 9616
rect 2834 9560 2839 9616
rect 0 9558 2839 9560
rect 0 9528 800 9558
rect 2773 9555 2839 9558
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 6637 778 6703 781
rect 7543 778 8343 808
rect 6637 776 8343 778
rect 6637 720 6642 776
rect 6698 720 8343 776
rect 6637 718 8343 720
rect 6637 715 6703 718
rect 7543 688 8343 718
<< via3 >>
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 8192 4528 8208
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 7648 5188 8208
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__clkbuf_2  _14_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3864 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _15_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 4692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _16_
timestamp 1693170804
transform 1 0 5888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _17_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 5428 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _18_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 5428 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o32ai_1  _19_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 4600 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _20_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _21_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _22_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 4600 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _23_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 4324 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _24_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _25_
timestamp 1693170804
transform 1 0 4968 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _26_
timestamp 1693170804
transform 1 0 3864 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor4b_1  _27_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 5428 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _28_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 5888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _29_
timestamp 1693170804
transform -1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _30_
timestamp 1693170804
transform -1 0 2576 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _31_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 2944 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_2  _32_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3956 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _33_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 1748 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _34_
timestamp 1693170804
transform 1 0 1472 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clock_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 2576 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1693170804
transform -1 0 6256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1693170804
transform -1 0 6716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 2760 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clock
timestamp 1693170804
transform -1 0 3312 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clock
timestamp 1693170804
transform 1 0 2760 0 -1 6528
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1693170804
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1693170804
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1693170804
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_61
timestamp 1693170804
transform 1 0 6716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_3
timestamp 1693170804
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_24
timestamp 1693170804
transform 1 0 3312 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_28
timestamp 1693170804
transform 1 0 3680 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_33 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 4140 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1693170804
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1693170804
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1693170804
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1693170804
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_15
timestamp 1693170804
transform 1 0 2484 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1693170804
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_29
timestamp 1693170804
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 4232 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_51
timestamp 1693170804
transform 1 0 5796 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_3
timestamp 1693170804
transform 1 0 1380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_24
timestamp 1693170804
transform 1 0 3312 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_35
timestamp 1693170804
transform 1 0 4324 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_45
timestamp 1693170804
transform 1 0 5244 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_53
timestamp 1693170804
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_57
timestamp 1693170804
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1693170804
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_15
timestamp 1693170804
transform 1 0 2484 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_18
timestamp 1693170804
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 1693170804
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_29
timestamp 1693170804
transform 1 0 3772 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_36
timestamp 1693170804
transform 1 0 4416 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_42
timestamp 1693170804
transform 1 0 4968 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_46
timestamp 1693170804
transform 1 0 5336 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_50
timestamp 1693170804
transform 1 0 5704 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_55
timestamp 1693170804
transform 1 0 6164 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_3
timestamp 1693170804
transform 1 0 1380 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_11
timestamp 1693170804
transform 1 0 2116 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_16
timestamp 1693170804
transform 1 0 2576 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_38
timestamp 1693170804
transform 1 0 4600 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_50
timestamp 1693170804
transform 1 0 5704 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_57
timestamp 1693170804
transform 1 0 6348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_3
timestamp 1693170804
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1693170804
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_29
timestamp 1693170804
transform 1 0 3772 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_33
timestamp 1693170804
transform 1 0 4140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_45
timestamp 1693170804
transform 1 0 5244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_57
timestamp 1693170804
transform 1 0 6348 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1693170804
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_15
timestamp 1693170804
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_38
timestamp 1693170804
transform 1 0 4600 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_47
timestamp 1693170804
transform 1 0 5428 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_52
timestamp 1693170804
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_57
timestamp 1693170804
transform 1 0 6348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_3
timestamp 1693170804
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_20
timestamp 1693170804
transform 1 0 2944 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_25
timestamp 1693170804
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_29
timestamp 1693170804
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_52
timestamp 1693170804
transform 1 0 5888 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_60
timestamp 1693170804
transform 1 0 6624 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1693170804
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1693170804
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1693170804
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1693170804
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1693170804
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1693170804
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_57
timestamp 1693170804
transform 1 0 6348 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_3
timestamp 1693170804
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_20
timestamp 1693170804
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1693170804
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1693170804
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_53
timestamp 1693170804
transform 1 0 5980 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_57
timestamp 1693170804
transform 1 0 6348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_62
timestamp 1693170804
transform 1 0 6808 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1693170804
transform -1 0 6808 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 6164 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_12  output3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 2944 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_11
timestamp 1693170804
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1693170804
transform -1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_12
timestamp 1693170804
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1693170804
transform -1 0 7176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_13
timestamp 1693170804
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1693170804
transform -1 0 7176 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_14
timestamp 1693170804
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1693170804
transform -1 0 7176 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_15
timestamp 1693170804
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1693170804
transform -1 0 7176 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_16
timestamp 1693170804
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1693170804
transform -1 0 7176 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_17
timestamp 1693170804
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1693170804
transform -1 0 7176 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_18
timestamp 1693170804
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1693170804
transform -1 0 7176 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_19
timestamp 1693170804
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1693170804
transform -1 0 7176 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_20
timestamp 1693170804
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1693170804
transform -1 0 7176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_21
timestamp 1693170804
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1693170804
transform -1 0 7176 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_23
timestamp 1693170804
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_24
timestamp 1693170804
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_25
timestamp 1693170804
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_26
timestamp 1693170804
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_27
timestamp 1693170804
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_28
timestamp 1693170804
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_29
timestamp 1693170804
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_30
timestamp 1693170804
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_31
timestamp 1693170804
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_32
timestamp 1693170804
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_33
timestamp 1693170804
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_34
timestamp 1693170804
transform 1 0 6256 0 1 7616
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 8208 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 8208 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 clock
port 2 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 detector_out
port 3 nsew signal tristate
flabel metal2 s 7746 9687 7802 10487 0 FreeSans 224 90 0 0 reset
port 4 nsew signal input
flabel metal3 s 7543 688 8343 808 0 FreeSans 480 0 0 0 sequence_in
port 5 nsew signal input
rlabel metal1 4140 7616 4140 7616 0 VGND
rlabel metal1 4140 8160 4140 8160 0 VPWR
rlabel metal1 5658 6426 5658 6426 0 _00_
rlabel metal1 3220 6630 3220 6630 0 _01_
rlabel metal2 2438 4590 2438 4590 0 _02_
rlabel metal1 2622 6392 2622 6392 0 _03_
rlabel metal2 4094 3196 4094 3196 0 _04_
rlabel metal1 4922 3978 4922 3978 0 _05_
rlabel metal1 5934 4114 5934 4114 0 _06_
rlabel metal2 5566 5508 5566 5508 0 _07_
rlabel metal1 4830 4114 4830 4114 0 _08_
rlabel metal1 3864 2890 3864 2890 0 _09_
rlabel metal1 4048 4250 4048 4250 0 _10_
rlabel metal1 3726 4012 3726 4012 0 _11_
rlabel metal1 4462 3978 4462 3978 0 _12_
rlabel metal1 4968 3706 4968 3706 0 _13_
rlabel metal1 3450 5338 3450 5338 0 clknet_0_clock
rlabel metal2 1518 4896 1518 4896 0 clknet_1_0__leaf_clock
rlabel metal1 4002 6732 4002 6732 0 clknet_1_1__leaf_clock
rlabel metal1 1334 4454 1334 4454 0 clock
rlabel metal1 4876 6222 4876 6222 0 current_state\[0\]
rlabel metal2 3542 6018 3542 6018 0 current_state\[1\]
rlabel metal1 3082 3638 3082 3638 0 current_state\[2\]
rlabel metal1 2507 7922 2507 7922 0 detector_out
rlabel metal1 2530 5236 2530 5236 0 net1
rlabel metal1 5750 3570 5750 3570 0 net2
rlabel metal2 2806 7242 2806 7242 0 net3
rlabel metal2 4738 5474 4738 5474 0 next_state\[0\]
rlabel metal1 3910 5780 3910 5780 0 next_state\[1\]
rlabel metal2 3358 4250 3358 4250 0 next_state\[2\]
rlabel metal1 7222 7854 7222 7854 0 reset
rlabel metal2 6670 1513 6670 1513 0 sequence_in
<< properties >>
string FIXED_BBOX 0 0 8343 10487
<< end >>
